module ALUSrcMUX();

endmodule

module ALUOp();

endmodule

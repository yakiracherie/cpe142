module PCAdder();

endmodule

module HazardDetection();

endmodule

module RegDstMUX.v();

endmodule

module PC();

endmodule

module BranchAND();

endmodule

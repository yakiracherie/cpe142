module BranchMUX();

endmodule

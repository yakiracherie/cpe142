module JumpMUX();

endmodule
